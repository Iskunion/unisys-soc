`ifndef _PERFS
`define _PERFS

//masters
`define CPU_NO 0

//slaves
`define MAINMEM_NO 0
`define UART_NO    1


`endif