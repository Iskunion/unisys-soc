`ifndef _TIMER
`define _TIMER

`include "uibi.sv"

module timer(
  input wire clk,
  input wire rst,
  `UIBI_SLAVE
);

endmodule

`endif