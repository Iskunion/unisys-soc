`ifndef _PERFS
`define _PERFS

`define CPU_NO 0

`endif