`ifndef _MAINMEM
`define _MAINMEM
`endif